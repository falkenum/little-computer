
`timescale 1us / 1ps

module i2c(
	input clk, 
	input [7:0] data_in,
	output scl,
	output [7:0] data_out,
	inout sda
	);

endmodule