
`include "defs.vh"

`timescale 1 ns / 1 ps
module lc_tb;
endmodule

